module pc_plus_4 (
    input   [31:0]  pc,
    output  [31:0]  pcplus4
);

assign pcplus4 = pc + 32'd4;

endmodule